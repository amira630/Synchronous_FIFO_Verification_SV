interface FIFO_if;
    
endinterface